//------------------------------------------------------------------------------
// SPDX-License-Identifier: GPL-3.0-or-later
// SPDX-FileType: SOURCE
// SPDX-FileCopyrightText: (c) 2022, antongale
//------------------------------------------------------------------------------

`default_nettype none

module slapfight ();

endmodule
